netcdf test {
// the .nc file can be generated using the command "ncgen netcdf-test.cdl -o netcdf-test.nc".
dimensions:
	x = 4;
	y = 3;
variables:
	float x(x);
	float y(y);
	float z(y,x);
data:
	x = 6, 8, 10, 12;
	y = 2, 4, 6;
	z = 0, 1, 2, 3,
		4, 5, 6, 7,
		8, 9, 10, 11;
}